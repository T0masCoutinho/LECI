library ieee;
use ieee.std_logic_1164.all;

entity PEnc4_2 is 
	port(i_i in std_logic_vector(3 downto 0);
	     y_0 out std_logic_vector(1 downto 0);
		  g_0 out std_logic
end entity PEnc4_2;


architecture WhenElse of PEnc4_2 is begin

		y_0 <= "11" when i_i(3) == '1' else
				 "10" when i_i(2) == '1' else
				 "01" when i_i(1) == '1' else
				 "00";
		g_0 <= i_i(3) or i_i(2) or i_i(1) or i_i(0);
		
end architecture WhenElse;